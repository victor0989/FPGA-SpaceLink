`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11.02.2025 05:53:07
// Design Name: 
// Module Name: disp_hex_mux
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module disp_hex_mux(
    input clk,
    input reset,
    input [3:0] hex3,
    input [3:0] hex2,
    input [3:0] hex1,
    input [3:0] hex0,
    input [3:0] dp_in,
    input [3:0] an,
    input [7:0] sseg
    );
endmodule
